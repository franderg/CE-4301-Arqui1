module sevenSeg(R,Seg);
	
	input [3:0] R;

	output reg [6:0] Seg;

	always @ (R)begin
		case (R)
			4'd0 :  Seg = 7'b1000000;
			4'd1 :  Seg = 7'b1111001;
			4'd2 :  Seg = 7'b0100100;
			4'd3 :  Seg = 7'b0110000;
			4'd4 :  Seg = 7'b0011001;
			4'd5 :  Seg = 7'b0010010;
			4'd6 :  Seg = 7'b0000010;
			4'd7 :  Seg = 7'b1111000;
			4'd8 :  Seg = 7'b0000000;
			4'd9 :  Seg = 7'b0010000;
			4'd10 :  Seg = 7'b0001000;
			4'd11 :  Seg = 7'b0000011;
			4'd12 :  Seg = 7'b1000110;
			4'd13 :  Seg = 7'b0100001;
			4'd14 :  Seg = 7'b0000110;
			4'd15 :  Seg = 7'b0001110;
			default :  Seg = 7'b1000000;
		endcase
	end
endmodule


//			4'b0000 :  Seg = 7b'0000001;
//			4'b0001 :  Seg = 7b'1001111;
//			4'b0010 :  Seg = 7b'0010010;
//			4'b0011 :  Seg = 7b'0000110;
//			4'b0100 :  Seg = 7b'1001100;
//			4'b0101 :  Seg = 7b'0100000;
//			4'b0111 :  Seg = 7b'0001111;
//			4'b1000 :  Seg = 7b'0000000;
//			4'b1001 :  Seg = 7b'0001100;
//			4'b1010 :  Seg = 7b'0001000;
//			4'b1011 :  Seg = 7b'1100000;
//			4'b1100 :  Seg = 7b'0000111;
//			4'b1101 :  Seg = 7b'1000010;
//			4'b1110 :  Seg = 7b'0011000;
//			4'b1111 :  Seg = 7b'0000000;
//			default :  Seg = 7b'1111111;