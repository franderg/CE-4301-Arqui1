// unsaved.v

// Generated using ACDS version 17.0 595

`timescale 1 ps / 1 ps
module unsaved (
		input  wire        clk_clk,         //   clk.clk
		input  wire [4:0]  pc_address,      //    pc.address
		input  wire        pc_debugaccess,  //      .debugaccess
		input  wire        pc_clken,        //      .clken
		input  wire        pc_chipselect,   //      .chipselect
		input  wire        pc_write,        //      .write
		output wire [31:0] pc_readdata,     //      .readdata
		input  wire [31:0] pc_writedata,    //      .writedata
		input  wire [3:0]  pc_byteenable,   //      .byteenable
		input  wire        reset_reset,     // reset.reset
		input  wire        reset_reset_req  //      .reset_req
	);

	unsaved_onchip_memory2_0 onchip_memory2_0 (
		.clk         (clk_clk),         //   clk1.clk
		.address     (pc_address),      //     s1.address
		.debugaccess (pc_debugaccess),  //       .debugaccess
		.clken       (pc_clken),        //       .clken
		.chipselect  (pc_chipselect),   //       .chipselect
		.write       (pc_write),        //       .write
		.readdata    (pc_readdata),     //       .readdata
		.writedata   (pc_writedata),    //       .writedata
		.byteenable  (pc_byteenable),   //       .byteenable
		.reset       (reset_reset),     // reset1.reset
		.reset_req   (reset_reset_req), //       .reset_req
		.freeze      (1'b0)             // (terminated)
	);

endmodule
