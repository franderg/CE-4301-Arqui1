module sevenSeg(R,Seg);
	
	input [3:0] R;

	output reg [6:0] Seg;

	always @ (R)begin
		case (R)
			4'b0000 :  Seg = 7'b1111110;
			4'b0001 :  Seg = 7'b0110000;
			4'b0010 :  Seg = 7'b1101101;
			4'b0011 :  Seg = 7'b1111001;
			4'b0100 :  Seg = 7'b0110011;
			4'b0101 :  Seg = 7'b1011011;
			4'b0110 :  Seg = 7'b1011111;
			4'b0111 :  Seg = 7'b1110000;
			4'b1000 :  Seg = 7'b1111111;
			4'b1001 :  Seg = 7'b1110011;
			4'b1010 :  Seg = 7'b1110111;
			4'b1011 :  Seg = 7'b0011111;
			4'b1100 :  Seg = 7'b1111000;
			4'b1101 :  Seg = 7'b1100111;
			4'b1111 :  Seg = 7'b1111111;
			default :  Seg = 7'b0000000;
		endcase
	end
endmodule



//			4'b0000 :  Seg = 7b'0000001;
//			4'b0001 :  Seg = 7b'1001111;
//			4'b0010 :  Seg = 7b'0010010;
//			4'b0011 :  Seg = 7b'0000110;
//			4'b0100 :  Seg = 7b'1001100;
//			4'b0101 :  Seg = 7b'0100000;
//			4'b0111 :  Seg = 7b'0001111;
//			4'b1000 :  Seg = 7b'0000000;
//			4'b1001 :  Seg = 7b'0001100;
//			4'b1010 :  Seg = 7b'0001000;
//			4'b1011 :  Seg = 7b'1100000;
//			4'b1100 :  Seg = 7b'0000111;
//			4'b1101 :  Seg = 7b'1000010;
//			4'b1110 :  Seg = 7b'0011000;
//			4'b1111 :  Seg = 7b'0000000;
//			default :  Seg = 7b'1111111;